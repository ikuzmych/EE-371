module binarySearch(); 


endmodule 



module binarySearch_testbench();




endmodule
